entity test is
end entity;

architecture rtl of test is
begin
end rtl;

architecture rtl2 of test is
begin
end rtl2;
