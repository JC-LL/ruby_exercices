entity test2 is
  port(
    reset_n : in bit;
    clk : in boolean;
    a,b : in bit
  );
end entity;

architecture rtl of test is
begin
end rtl;
